    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   Saver+Position   xyz      t���r��  ��